use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.tcp_common.all;

entity application is
  port(
       clk : in std_ulogic;
	   reset: in std_ulogic;
	   
       o_start          :  out std_ulogic;
	   o_active_mode  :  out  std_ulogic;
	   o_open         :  out std_ulogic;     
	   o_timeout      :  out  unsigned (10 downto 0);
	   i_close        :  in  std_ulogic;
	   ---------------------------------------------
	   -- SRC IP,PORT / DST IP,PORT defined by App 
	   ---------------------------------------------
	   o_src_ip       : out   t_ipv4_address;
	   o_dst_ip       : out   t_ipv4_address;
	   o_src_port     : out   t_tcp_port;
	   o_dst_port     : out   t_tcp_port;
	   
       rx_tdata: in std_ulogic_vector(7 downto 0);
       rx_tvalid: in std_ulogic;
	   rx_tready: out std_ulogic;
	   rx_tlast: in std_ulogic;
	   
	   tx_tdata: out std_ulogic_vector(7 downto 0);
	   tx_tvalid: out std_ulogic;
	   tx_tready: in std_ulogic;
	   tx_tlast: out std_ulogic
	   );
	   
end application;

architecture behavioural of application is

type FRAME1 is array(0 to 50) of std_ulogic_vector(7 downto 0);
type FRAME2 is array(0 to 4200) of std_ulogic_vector(7 downto 0);
type FRAME3 is array(0 to 1400) of std_ulogic_vector(7 downto 0);

type state_t is (start_trans, send_frame1, send_frame2, send_frame3, request_close);
signal state: state_t;
signal i: integer:= 0;

signal frame_1: FRAME1 := (X"12", X"DC", X"17", X"BC", X"B7", X"5D", X"58", X"72", X"59", X"A0", X"0F", X"33", X"35", X"B9", X"BA", X"5B", X"D8", X"82", X"FD", X"3A", X"FD", X"51", X"64", X"47", X"37", X"35", X"24", X"CE", X"1E", X"B6", X"76", X"95", X"6B", X"6E", X"3C", X"96", X"72", X"37", X"95", X"A2", X"3A", X"8D", X"86", X"B3", X"F7", X"28", X"28", X"D4", X"7E", X"7B", X"95");
signal frame_2: FRAME2 := (X"51", X"EC", X"3C", X"33", X"E7", X"C5", X"F4", X"99", X"4E", X"19", X"6A", X"B8", X"12", X"03", X"E2", X"7C", X"7A", X"8E", X"F5", X"BD", X"B4", X"87", X"78", X"A3", X"05", X"27", X"6A", X"13", X"79", X"A6", X"0A", X"F9", X"53", X"67", X"81", X"99", X"3B", X"CF", X"3C", X"D3", X"59", X"93", X"2E", X"60", X"6A", X"11", X"C7", X"B6", X"D3", X"D8", X"33", X"B4", X"E6", X"15", X"57", X"02", X"13", X"AF", X"C6", X"69", X"20", X"C1", X"54", X"99", X"EA", X"34", X"8A", X"0A", X"7E", X"35", X"42", X"36", X"BC", X"FD", X"B6", X"28", X"BD", X"FD", X"4E", X"7E", X"85", X"46", X"B6", X"E2", X"B7", X"8A", X"77", X"50", X"58", X"2C", X"7E", X"5D", X"C7", X"29", X"38", X"01", X"71", X"D4", X"4B", X"AC", X"75", X"1B", X"25", X"43", X"E1", X"5B", X"59", X"FE", X"FC", X"A1", X"E9", X"5F", X"F1", X"10", X"3D", X"98", X"18", X"22", X"DE", X"D7", X"0C", X"06", X"1D", X"6F", X"44", X"F8", X"E7", X"9C", X"FC", X"D6", X"AC", X"AD", X"DE", X"FE", X"F7", X"BD", X"17", X"EE", X"E5", X"FE", X"EB", X"EC", X"60", X"63", X"9A", X"52", X"96", X"2C", X"51", X"9C", X"65", X"65", X"7A", X"0E", X"52", X"15", X"BA", X"DB", X"2F", X"69", X"C6", X"6A", X"0A", X"AA", X"8D", X"8C", X"0F", X"A2", X"83", X"20", X"A7", X"A7", X"91", X"7F", X"B9", X"CD", X"3D", X"72", X"D0", X"C1", X"B2", X"D1", X"4F", X"F9", X"02", X"5E", X"87", X"D0", X"73", X"C6", X"2F", X"7F", X"97", X"6D", X"EC", X"65", X"61", X"3F", X"88", X"49", X"02", X"8D", X"75", X"70", X"48", X"27", X"67", X"25", X"13", X"E8", X"63", X"55", X"5B", X"06", X"D1", X"1F", X"2F", X"F7", X"88", X"E5", X"89", X"61", X"4A", X"25", X"81", X"50", X"A5", X"3A", X"B3", X"9C", X"73", X"D8", X"62", X"1D", X"63", X"9E", X"C6", X"CF", X"1A", X"BE", X"A8", X"FB", X"A7", X"35", X"53", X"4E", X"8B", X"B7", X"A5", X"2C", X"DB", X"B5", X"EC", X"8A", X"5E", X"B3", X"D1", X"8A", X"5D", X"9D", X"B9", X"75", X"CE", X"E3", X"97", X"BD", X"57", X"F9", X"E1", X"EE", X"20", X"CA", X"23", X"15", X"B0", X"50", X"41", X"21", X"F6", X"57", X"36", X"60", X"F6", X"31", X"8B", X"AE", X"31", X"9E", X"E5", X"10", X"B2", X"CB", X"C9", X"7E", X"40", X"FE", X"FE", X"62", X"F2", X"B4", X"C3", X"7A", X"5B", X"2B", X"75", X"73", X"F3", X"42", X"A6", X"42", X"12", X"3A", X"A3", X"58", X"3B", X"84", X"1D", X"AC", X"94", X"69", X"25", X"7F", X"9B", X"A1", X"57", X"5D", X"A0", X"56", X"1C", X"4F", X"F2", X"C5", X"11", X"D1", X"6C", X"E7", X"CB", X"10", X"64", X"99", X"40", X"12", X"66", X"69", X"85", X"62", X"99", X"C4", X"F3", X"D9", X"93", X"C6", X"DC", X"A7", X"BF", X"8D", X"A2", X"D3", X"1D", X"7F", X"73", X"18", X"4E", X"5E", X"62", X"17", X"BF", X"9E", X"FB", X"43", X"3E", X"60", X"FF", X"DF", X"B7", X"D6", X"41", X"A0", X"12", X"60", X"3B", X"E3", X"81", X"04", X"37", X"2B", X"42", X"1B", X"AD", X"CE", X"5D", X"4C", X"EC", X"0D", X"9E", X"84", X"52", X"21", X"3B", X"7E", X"8D", X"4D", X"11", X"3A", X"05", X"E3", X"73", X"9A", X"5E", X"D8", X"2C", X"0D", X"56", X"B9", X"D4", X"D2", X"B9", X"CD", X"02", X"69", X"1A", X"68", X"71", X"06", X"A1", X"05", X"34", X"48", X"AA", X"18", X"F7", X"93", X"C2", X"67", X"3D", X"11", X"1A", X"13", X"EE", X"0F", X"8D", X"23", X"0D", X"6F", X"38", X"E2", X"20", X"82", X"0A", X"AC", X"47", X"15", X"13", X"4D", X"6D", X"41", X"64", X"D0", X"DF", X"B6", X"48", X"80", X"8E", X"77", X"6A", X"A2", X"FA", X"BA", X"1B", X"6D", X"0A", X"3D", X"B9", X"82", X"53", X"D2", X"74", X"E5", X"23", X"6F", X"C4", X"9D", X"08", X"C1", X"52", X"6C", X"63", X"A4", X"32", X"DA", X"F7", X"D2", X"8B", X"77", X"0E", X"FD", X"A7", X"FA", X"1C", X"15", X"0D", X"70", X"EC", X"ED", X"BF", X"7E", X"42", X"66", X"12", X"39", X"46", X"7B", X"7B", X"0F", X"1C", X"37", X"DC", X"E1", X"F5", X"17", X"33", X"42", X"B4", X"6B", X"65", X"90", X"F4", X"1A", X"11", X"AA", X"31", X"8B", X"ED", X"02", X"D5", X"E2", X"2C", X"24", X"F5", X"57", X"CD", X"90", X"C6", X"4D", X"E6", X"2C", X"E7", X"CD", X"84", X"8E", X"A7", X"BE", X"D3", X"CA", X"DB", X"7E", X"A5", X"F6", X"1B", X"F4", X"DD", X"26", X"BF", X"B4", X"A0", X"CB", X"59", X"43", X"62", X"B9", X"E8", X"D1", X"07", X"24", X"67", X"44", X"C9", X"FC", X"5D", X"39", X"82", X"7C", X"C5", X"2F", X"64", X"B0", X"CD", X"0C", X"16", X"B5", X"F4", X"13", X"B5", X"2E", X"1E", X"2C", X"3D", X"33", X"57", X"8B", X"7A", X"F4", X"AB", X"06", X"0B", X"E4", X"93", X"27", X"96", X"A7", X"90", X"EE", X"41", X"F5", X"9D", X"ED", X"90", X"D7", X"DB", X"69", X"86", X"ED", X"8F", X"9E", X"8B", X"99", X"F2", X"89", X"F3", X"09", X"ED", X"86", X"13", X"C6", X"8E", X"B7", X"17", X"91", X"E4", X"66", X"8A", X"41", X"4A", X"9E", X"26", X"25", X"27", X"6C", X"CF", X"7D", X"9F", X"A9", X"76", X"49", X"09", X"46", X"FF", X"87", X"C3", X"BB", X"85", X"B0", X"45", X"13", X"64", X"FB", X"FD", X"D0", X"1C", X"A8", X"8F", X"4D", X"D8", X"ED", X"D7", X"17", X"0F", X"E2", X"6B", X"57", X"46", X"BC", X"EA", X"37", X"FB", X"A9", X"13", X"BF", X"DD", X"44", X"B3", X"A9", X"37", X"DD", X"B6", X"66", X"38", X"3F", X"DE", X"FE", X"2F", X"68", X"14", X"62", X"43", X"31", X"23", X"B0", X"8E", X"6C", X"A2", X"50", X"3F", X"9A", X"4F", X"06", X"4B", X"B7", X"91", X"E9", X"88", X"C3", X"6E", X"6F", X"4F", X"C7", X"9D", X"2A", X"8E", X"CA", X"CC", X"B6", X"7B", X"3D", X"5F", X"B1", X"CF", X"80", X"44", X"2B", X"76", X"FB", X"7D", X"73", X"C3", X"95", X"69", X"6C", X"2D", X"D0", X"D1", X"4C", X"47", X"73", X"DE", X"1F", X"7B", X"A4", X"C6", X"F7", X"5B", X"6F", X"0B", X"8E", X"4F", X"32", X"7B", X"51", X"D8", X"7E", X"62", X"5A", X"75", X"CB", X"96", X"6D", X"3A", X"C5", X"99", X"B4", X"F5", X"9C", X"F8", X"61", X"B1", X"E4", X"B2", X"1D", X"23", X"31", X"BB", X"D4", X"8C", X"6F", X"CA", X"9F", X"0B", X"05", X"16", X"27", X"7D", X"58", X"AD", X"8A", X"29", X"72", X"A7", X"FC", X"34", X"1E", X"86", X"19", X"BD", X"91", X"59", X"A9", X"FB", X"63", X"70", X"13", X"CB", X"F1", X"DF", X"37", X"06", X"6F", X"1F", X"8C", X"CE", X"73", X"14", X"1C", X"C9", X"5E", X"15", X"FF", X"5A", X"FE", X"E1", X"42", X"59", X"FB", X"A3", X"8D", X"6B", X"4F", X"87", X"45", X"27", X"65", X"88", X"AE", X"40", X"C9", X"D0", X"D6", X"A4", X"06", X"AB", X"FA", X"52", X"6D", X"4C", X"9F", X"0B", X"39", X"31", X"12", X"70", X"F4", X"DD", X"37", X"FB", X"7C", X"19", X"DE", X"5F", X"8A", X"3A", X"49", X"63", X"58", X"4C", X"76", X"99", X"14", X"A2", X"E1", X"BE", X"5B", X"C8", X"B6", X"FF", X"77", X"13", X"F9", X"D8", X"8C", X"E4", X"FB", X"FD", X"2A", X"27", X"73", X"54", X"E1", X"B1", X"C5", X"D1", X"ED", X"A9", X"1E", X"B0", X"01", X"62", X"16", X"3A", X"FB", X"B4", X"4F", X"7A", X"20", X"A9", X"8B", X"17", X"EC", X"CE", X"67", X"76", X"97", X"EA", X"DD", X"A1", X"B9", X"FA", X"98", X"37", X"BF", X"93", X"00", X"9D", X"95", X"A1", X"23", X"B1", X"37", X"73", X"1E", X"F9", X"E1", X"ED", X"15", X"CB", X"41", X"CA", X"67", X"9E", X"57", X"A0", X"7F", X"1A", X"9C", X"98", X"1C", X"8C", X"71", X"50", X"B1", X"7F", X"13", X"82", X"5D", X"3A", X"AE", X"22", X"35", X"E4", X"BC", X"D8", X"88", X"1A", X"A5", X"60", X"80", X"4B", X"E9", X"3B", X"0A", X"1A", X"DC", X"DC", X"D9", X"51", X"1F", X"A2", X"46", X"E3", X"4F", X"D2", X"D9", X"F6", X"2C", X"D3", X"A4", X"14", X"9F", X"C1", X"27", X"5F", X"A5", X"4F", X"DE", X"7D", X"ED", X"96", X"74", X"96", X"14", X"19", X"F9", X"BC", X"6B", X"32", X"A2", X"F7", X"99", X"FA", X"5A", X"81", X"A7", X"7D", X"C0", X"8C", X"B5", X"EE", X"90", X"4D", X"DA", X"26", X"DA", X"60", X"E3", X"E5", X"77", X"88", X"F2", X"C9", X"E0", X"3C", X"B4", X"CF", X"5E", X"42", X"4B", X"60", X"EA", X"66", X"BA", X"8B", X"BB", X"DA", X"13", X"F3", X"74", X"33", X"76", X"FE", X"76", X"A2", X"EA", X"DE", X"BB", X"DE", X"73", X"52", X"AA", X"C2", X"A0", X"45", X"03", X"91", X"74", X"3D", X"4B", X"CF", X"30", X"BA", X"E7", X"6C", X"5A", X"13", X"C2", X"B3", X"81", X"28", X"17", X"6F", X"00", X"64", X"DF", X"DC", X"0D", X"A8", X"BE", X"3B", X"6D", X"84", X"31", X"86", X"A9", X"AB", X"07", X"13", X"27", X"B9", X"9E", X"35", X"6A", X"93", X"7A", X"88", X"02", X"F6", X"C6", X"BF", X"42", X"FE", X"4C", X"C8", X"28", X"CA", X"8A", X"69", X"B2", X"F4", X"BB", X"3E", X"16", X"28", X"30", X"35", X"65", X"BB", X"6C", X"BE", X"56", X"D8", X"A3", X"EA", X"AB", X"C5", X"39", X"36", X"39", X"C8", X"F8", X"BC", X"65", X"55", X"D6", X"6D", X"97", X"3A", X"EB", X"3D", X"95", X"ED", X"A1", X"A2", X"62", X"75", X"53", X"06", X"18", X"A5", X"38", X"E0", X"29", X"87", X"DE", X"60", X"9F", X"AA", X"3F", X"16", X"70", X"FF", X"0A", X"B1", X"1D", X"71", X"D9", X"C2", X"6C", X"28", X"CD", X"24", X"47", X"12", X"8B", X"08", X"68", X"86", X"C9", X"EC", X"16", X"D7", X"3F", X"8B", X"24", X"55", X"33", X"53", X"92", X"12", X"86", X"37", X"CB", X"7B", X"DD", X"8D", X"65", X"77", X"40", X"57", X"D1", X"65", X"0F", X"51", X"3B", X"8D", X"4D", X"16", X"FE", X"4D", X"33", X"DC", X"28", X"7B", X"81", X"7D", X"47", X"50", X"9F", X"11", X"62", X"50", X"39", X"C3", X"D9", X"C5", X"A6", X"D6", X"A5", X"12", X"5D", X"31", X"E5", X"2D", X"F9", X"77", X"73", X"E2", X"9A", X"61", X"FF", X"B2", X"B8", X"A8", X"CE", X"CA", X"84", X"D9", X"68", X"CA", X"B0", X"E9", X"12", X"58", X"08", X"7E", X"BA", X"DB", X"C0", X"EC", X"3D", X"80", X"41", X"2F", X"A7", X"F1", X"0E", X"75", X"68", X"3F", X"C9", X"2E", X"CC", X"A7", X"1E", X"0D", X"30", X"F5", X"3F", X"50", X"CA", X"3B", X"EF", X"8E", X"93", X"08", X"4A", X"54", X"BB", X"04", X"66", X"0D", X"EA", X"0F", X"61", X"8C", X"7F", X"74", X"F7", X"DF", X"A4", X"83", X"23", X"CE", X"8B", X"02", X"55", X"6C", X"87", X"36", X"AB", X"A1", X"5F", X"31", X"65", X"78", X"0C", X"AC", X"E5", X"65", X"6C", X"49", X"DC", X"60", X"9E", X"3E", X"EC", X"77", X"7C", X"A7", X"3F", X"B1", X"DD", X"2E", X"73", X"E7", X"10", X"BE", X"A9", X"28", X"43", X"84", X"9D", X"FB", X"25", X"E9", X"80", X"B4", X"5B", X"5C", X"BA", X"CC", X"50", X"85", X"07", X"8C", X"C8", X"A9", X"D8", X"AE", X"91", X"A5", X"6B", X"23", X"9A", X"45", X"B3", X"E7", X"1C", X"71", X"76", X"21", X"4A", X"D8", X"AB", X"9D", X"7C", X"FD", X"3E", X"6F", X"B2", X"8F", X"1B", X"59", X"BB", X"F0", X"65", X"20", X"44", X"DB", X"37", X"6B", X"99", X"34", X"D1", X"D4", X"00", X"EB", X"76", X"FE", X"4A", X"98", X"D9", X"EE", X"89", X"77", X"9C", X"1F", X"CD", X"48", X"25", X"2A", X"35", X"01", X"44", X"C2", X"19", X"34", X"A4", X"D6", X"68", X"51", X"15", X"A0", X"73", X"D1", X"20", X"EC", X"58", X"C1", X"D7", X"AF", X"0C", X"C1", X"2F", X"FD", X"CF", X"2A", X"DC", X"56", X"9F", X"49", X"46", X"5A", X"39", X"24", X"FE", X"8F", X"33", X"C3", X"AE", X"28", X"B8", X"13", X"61", X"C3", X"A6", X"08", X"7B", X"95", X"F6", X"6E", X"F6", X"F7", X"58", X"24", X"61", X"BC", X"C7", X"37", X"99", X"18", X"85", X"8A", X"F9", X"C6", X"32", X"00", X"D6", X"83", X"A8", X"3B", X"EB", X"AD", X"67", X"5B", X"D1", X"14", X"1A", X"EE", X"20", X"4B", X"E3", X"16", X"4E", X"36", X"CF", X"A2", X"7F", X"EF", X"06", X"0C", X"0E", X"B7", X"36", X"5A", X"D1", X"C2", X"E2", X"55", X"A8", X"61", X"A3", X"DE", X"67", X"BC", X"5F", X"98", X"DD", X"AD", X"D8", X"B8", X"B8", X"73", X"92", X"01", X"A2", X"A3", X"2A", X"8D", X"58", X"A9", X"26", X"94", X"E0", X"2D", X"37", X"28", X"04", X"A4", X"1D", X"EB", X"FD", X"62", X"52", X"62", X"C0", X"23", X"AC", X"45", X"5D", X"BA", X"D2", X"B8", X"0E", X"4C", X"76", X"3F", X"3C", X"C6", X"1A", X"95", X"29", X"93", X"F2", X"93", X"F4", X"06", X"E3", X"74", X"35", X"9A", X"8E", X"47", X"F6", X"26", X"32", X"29", X"EA", X"07", X"A8", X"36", X"3A", X"6C", X"10", X"B7", X"6A", X"18", X"41", X"40", X"B0", X"77", X"C4", X"11", X"44", X"2F", X"74", X"B7", X"2A", X"B3", X"D7", X"5E", X"67", X"6B", X"55", X"A1", X"9E", X"E8", X"1C", X"84", X"73", X"E4", X"B5", X"35", X"A1", X"64", X"27", X"68", X"E2", X"C6", X"2B", X"5D", X"5A", X"03", X"6E", X"47", X"97", X"39", X"FF", X"E9", X"5C", X"CE", X"5C", X"87", X"81", X"5F", X"44", X"2F", X"24", X"8E", X"79", X"94", X"96", X"EF", X"89", X"E9", X"E7", X"B6", X"B2", X"79", X"15", X"A5", X"FC", X"8E", X"C3", X"81", X"3F", X"05", X"33", X"63", X"F1", X"53", X"CF", X"15", X"AD", X"48", X"57", X"52", X"38", X"8E", X"30", X"6F", X"6E", X"61", X"E4", X"46", X"68", X"02", X"9B", X"DE", X"DE", X"62", X"67", X"5B", X"87", X"18", X"10", X"86", X"74", X"47", X"77", X"20", X"DF", X"9E", X"77", X"DE", X"15", X"9B", X"41", X"3F", X"8A", X"94", X"7B", X"20", X"9B", X"29", X"46", X"04", X"50", X"34", X"EA", X"BE", X"07", X"DD", X"39", X"96", X"0C", X"93", X"03", X"ED", X"5D", X"B4", X"0D", X"AE", X"AD", X"A5", X"E5", X"E0", X"F0", X"22", X"B6", X"CF", X"99", X"62", X"A4", X"72", X"4C", X"8F", X"69", X"43", X"6F", X"92", X"03", X"0A", X"50", X"77", X"B6", X"85", X"B7", X"89", X"47", X"20", X"1B", X"32", X"05", X"23", X"6D", X"2A", X"54", X"02", X"D0", X"86", X"87", X"8E", X"42", X"5A", X"15", X"74", X"41", X"0B", X"D1", X"17", X"9A", X"A2", X"45", X"A9", X"1F", X"93", X"AD", X"E0", X"D2", X"0B", X"25", X"39", X"7E", X"A1", X"D0", X"A1", X"53", X"B3", X"18", X"A3", X"9A", X"E3", X"52", X"0F", X"45", X"D4", X"B0", X"F7", X"47", X"3D", X"25", X"E3", X"D0", X"C1", X"63", X"B3", X"38", X"A8", X"A7", X"43", X"D1", X"27", X"F9", X"07", X"83", X"ED", X"B0", X"E1", X"D8", X"5A", X"11", X"8B", X"0A", X"08", X"DD", X"96", X"15", X"3D", X"73", X"A8", X"49", X"37", X"B9", X"95", X"78", X"12", X"FE", X"4B", X"95", X"3E", X"CA", X"20", X"D0", X"EB", X"56", X"F9", X"3C", X"17", X"4C", X"A3", X"8D", X"C7", X"21", X"D1", X"82", X"91", X"50", X"94", X"38", X"E9", X"3A", X"40", X"6D", X"F1", X"9B", X"92", X"7A", X"7C", X"FA", X"12", X"C6", X"C9", X"7C", X"D4", X"99", X"5F", X"71", X"0B", X"B4", X"1D", X"4C", X"20", X"8B", X"E0", X"BF", X"93", X"4B", X"91", X"82", X"2A", X"8A", X"FC", X"36", X"5B", X"C7", X"5A", X"A2", X"C1", X"B8", X"BC", X"DC", X"E3", X"E0", X"97", X"2B", X"6D", X"B2", X"37", X"80", X"E1", X"A1", X"B8", X"A8", X"3E", X"84", X"BD", X"17", X"F1", X"CD", X"38", X"EC", X"17", X"54", X"4E", X"41", X"9A", X"DA", X"43", X"C3", X"02", X"E6", X"10", X"9D", X"C3", X"30", X"86", X"D8", X"22", X"DA", X"B9", X"9C", X"01", X"C2", X"A1", X"D1", X"FD", X"11", X"26", X"38", X"00", X"91", X"2A", X"B0", X"24", X"61", X"31", X"53", X"6D", X"D2", X"8C", X"95", X"2A", X"DD", X"5F", X"93", X"84", X"BA", X"DD", X"E0", X"31", X"98", X"C0", X"C8", X"0A", X"38", X"67", X"53", X"7E", X"8A", X"34", X"87", X"CA", X"61", X"CF", X"15", X"54", X"C5", X"72", X"E5", X"5D", X"D5", X"2D", X"88", X"60", X"60", X"92", X"9A", X"D2", X"3F", X"05", X"DC", X"9C", X"52", X"89", X"6E", X"C8", X"85", X"30", X"1D", X"22", X"AE", X"5E", X"CC", X"C9", X"25", X"A4", X"90", X"0C", X"87", X"E2", X"66", X"35", X"68", X"24", X"60", X"EC", X"D9", X"AC", X"40", X"63", X"6B", X"D3", X"B3", X"B6", X"DD", X"76", X"F3", X"25", X"4E", X"DE", X"22", X"44", X"23", X"85", X"3C", X"67", X"B5", X"49", X"4C", X"A0", X"D9", X"33", X"2A", X"98", X"80", X"44", X"B4", X"3F", X"B5", X"91", X"EE", X"82", X"BD", X"D4", X"26", X"47", X"6C", X"1E", X"9E", X"C4", X"2F", X"B8", X"C9", X"5B", X"84", X"9F", X"6E", X"3D", X"56", X"D1", X"99", X"EA", X"F3", X"7A", X"0C", X"08", X"C8", X"2A", X"D4", X"96", X"DD", X"11", X"59", X"9D", X"44", X"70", X"F1", X"61", X"FC", X"60", X"2D", X"92", X"A8", X"2C", X"64", X"82", X"BD", X"51", X"FF", X"DF", X"9A", X"8B", X"F3", X"DE", X"60", X"EC", X"7C", X"85", X"4D", X"98", X"35", X"06", X"84", X"4C", X"CD", X"27", X"01", X"BA", X"B4", X"A0", X"3D", X"14", X"05", X"C3", X"F2", X"EA", X"7D", X"86", X"98", X"4D", X"4F", X"72", X"82", X"71", X"25", X"D5", X"07", X"0B", X"DF", X"0F", X"DA", X"BE", X"0B", X"D9", X"E4", X"87", X"00", X"33", X"30", X"E1", X"79", X"38", X"7F", X"90", X"BD", X"FA", X"CA", X"FD", X"35", X"8E", X"0B", X"CD", X"0C", X"6B", X"D8", X"D6", X"AF", X"FA", X"44", X"8B", X"B6", X"0E", X"20", X"BE", X"9E", X"6E", X"13", X"9E", X"78", X"10", X"E3", X"67", X"FC", X"5A", X"CA", X"3E", X"8E", X"CC", X"F1", X"87", X"9E", X"7F", X"62", X"B4", X"41", X"F9", X"53", X"1B", X"FF", X"B4", X"23", X"AF", X"72", X"53", X"5E", X"A3", X"56", X"1B", X"19", X"CF", X"B9", X"EF", X"FE", X"C3", X"25", X"2B", X"B1", X"C8", X"58", X"9F", X"E7", X"1B", X"68", X"FD", X"5B", X"CD", X"F6", X"23", X"31", X"DD", X"2E", X"94", X"A1", X"46", X"1F", X"FA", X"BD", X"89", X"72", X"A2", X"69", X"40", X"58", X"F2", X"89", X"B1", X"7D", X"F5", X"9F", X"E7", X"2F", X"B1", X"E1", X"D2", X"D4", X"71", X"A9", X"08", X"03", X"FB", X"36", X"5F", X"46", X"11", X"6D", X"DC", X"0F", X"F3", X"0C", X"1A", X"BB", X"20", X"94", X"DC", X"85", X"52", X"56", X"31", X"11", X"47", X"A4", X"2C", X"97", X"9A", X"26", X"11", X"D2", X"C7", X"E4", X"FE", X"1C", X"8B", X"D9", X"0B", X"53", X"BC", X"2B", X"80", X"6E", X"76", X"BB", X"98", X"48", X"B1", X"F8", X"A4", X"EC", X"A6", X"38", X"D5", X"87", X"0B", X"4E", X"BC", X"E4", X"40", X"73", X"12", X"F5", X"4F", X"AA", X"BC", X"86", X"07", X"63", X"15", X"73", X"EA", X"3F", X"1A", X"C0", X"44", X"7F", X"67", X"94", X"9F", X"B6", X"56", X"BC", X"E5", X"93", X"D4", X"3E", X"44", X"CC", X"D9", X"D7", X"16", X"EE", X"53", X"C1", X"D3", X"A9", X"38", X"3C", X"E1", X"17", X"88", X"A2", X"48", X"11", X"F3", X"09", X"CC", X"10", X"53", X"57", X"07", X"B8", X"23", X"EE", X"00", X"55", X"81", X"7F", X"82", X"29", X"A0", X"4F", X"9F", X"40", X"24", X"83", X"49", X"A4", X"4F", X"07", X"6E", X"16", X"9C", X"F7", X"06", X"5D", X"CA", X"B1", X"54", X"19", X"3F", X"97", X"43", X"11", X"F1", X"55", X"41", X"AA", X"1C", X"C8", X"9E", X"6C", X"7F", X"40", X"AF", X"AB", X"2C", X"03", X"14", X"C9", X"34", X"D1", X"8C", X"7E", X"73", X"8D", X"6A", X"2C", X"32", X"2D", X"ED", X"5C", X"9F", X"CE", X"F7", X"8E", X"17", X"B4", X"69", X"BD", X"E1", X"8E", X"75", X"AE", X"E3", X"B9", X"3C", X"DB", X"CB", X"DF", X"06", X"F5", X"78", X"67", X"9F", X"6E", X"20", X"7D", X"91", X"A1", X"D1", X"C6", X"71", X"EB", X"2D", X"C6", X"EC", X"7D", X"53", X"21", X"A1", X"83", X"FC", X"D8", X"87", X"AB", X"A2", X"49", X"45", X"AF", X"E8", X"1B", X"BB", X"85", X"70", X"78", X"DB", X"0E", X"3B", X"0C", X"E3", X"EC", X"02", X"82", X"B3", X"66", X"2E", X"63", X"4A", X"0A", X"38", X"01", X"67", X"E8", X"24", X"40", X"34", X"9C", X"48", X"CC", X"22", X"7C", X"CA", X"5F", X"FB", X"CF", X"F4", X"1D", X"5D", X"2F", X"DA", X"73", X"14", X"44", X"8A", X"13", X"D4", X"17", X"A4", X"3D", X"37", X"6C", X"40", X"BC", X"D1", X"FB", X"6E", X"6D", X"46", X"9F", X"C2", X"84", X"AC", X"8F", X"97", X"34", X"82", X"30", X"82", X"B9", X"62", X"4D", X"A7", X"03", X"6D", X"5F", X"55", X"F8", X"94", X"0C", X"F6", X"9B", X"B4", X"1D", X"21", X"AA", X"D8", X"24", X"8C", X"7D", X"64", X"34", X"95", X"42", X"DC", X"D0", X"93", X"64", X"AE", X"E8", X"11", X"93", X"3E", X"C6", X"53", X"0B", X"43", X"BA", X"59", X"F5", X"15", X"BE", X"2A", X"26", X"47", X"87", X"A0", X"0E", X"11", X"C3", X"48", X"04", X"BE", X"0D", X"0A", X"CD", X"C8", X"08", X"31", X"D6", X"B3", X"44", X"B7", X"05", X"EC", X"87", X"98", X"DC", X"2A", X"5F", X"20", X"C2", X"D0", X"79", X"43", X"FA", X"3D", X"D9", X"A4", X"34", X"B6", X"D2", X"5E", X"32", X"6E", X"56", X"6F", X"44", X"FC", X"C2", X"AF", X"0B", X"7B", X"E1", X"F6", X"04", X"DF", X"20", X"90", X"19", X"63", X"00", X"E5", X"65", X"87", X"39", X"BC", X"DF", X"5C", X"5E", X"C1", X"0B", X"21", X"09", X"E0", X"A3", X"E9", X"36", X"CF", X"63", X"CE", X"B3", X"BC", X"93", X"F4", X"52", X"7C", X"C1", X"DB", X"D2", X"50", X"A7", X"D1", X"21", X"76", X"66", X"88", X"96", X"49", X"7E", X"C3", X"D2", X"B3", X"A1", X"42", X"26", X"61", X"BD", X"85", X"BA", X"76", X"7C", X"27", X"31", X"B0", X"12", X"F6", X"2B", X"3E", X"EF", X"4A", X"8F", X"74", X"7E", X"95", X"C7", X"8F", X"2A", X"4B", X"89", X"67", X"8F", X"B4", X"9E", X"73", X"48", X"AE", X"5D", X"0F", X"0A", X"41", X"F0", X"A9", X"8E", X"9A", X"56", X"54", X"9B", X"0C", X"6E", X"90", X"69", X"FB", X"6F", X"88", X"3C", X"43", X"FD", X"C9", X"DA", X"44", X"FD", X"EB", X"B1", X"BA", X"27", X"9D", X"CD", X"14", X"83", X"C1", X"A1", X"3A", X"73", X"AF", X"31", X"59", X"8C", X"30", X"CE", X"43", X"D3", X"F0", X"AA", X"51", X"F2", X"B9", X"C3", X"87", X"9E", X"8F", X"DE", X"BA", X"41", X"50", X"26", X"79", X"74", X"FA", X"E1", X"1C", X"0C", X"97", X"68", X"E3", X"D8", X"9C", X"23", X"AA", X"4A", X"06", X"C1", X"FF", X"11", X"A3", X"6B", X"AD", X"5E", X"99", X"34", X"3E", X"7B", X"A3", X"F9", X"A5", X"62", X"18", X"F0", X"0A", X"69", X"32", X"D5", X"CC", X"EA", X"B8", X"9E", X"4C", X"8C", X"F3", X"DB", X"2C", X"E2", X"2A", X"5E", X"4D", X"51", X"34", X"EB", X"48", X"F3", X"02", X"3B", X"A2", X"86", X"E3", X"FF", X"96", X"5D", X"D9", X"55", X"22", X"68", X"10", X"1B", X"22", X"D0", X"93", X"3E", X"47", X"C2", X"13", X"87", X"E3", X"AF", X"6D", X"97", X"62", X"8F", X"6C", X"14", X"CA", X"97", X"E8", X"8F", X"73", X"19", X"72", X"08", X"47", X"BA", X"F8", X"47", X"FA", X"ED", X"73", X"FB", X"18", X"93", X"C9", X"46", X"70", X"0C", X"82", X"2E", X"A9", X"98", X"52", X"6C", X"28", X"44", X"57", X"50", X"6F", X"C5", X"02", X"51", X"1C", X"F0", X"F2", X"1E", X"ED", X"73", X"F2", X"41", X"8E", X"B4", X"1D", X"7D", X"F6", X"59", X"78", X"50", X"8B", X"F5", X"51", X"8E", X"AE", X"05", X"32", X"71", X"11", X"94", X"43", X"87", X"AF", X"01", X"68", X"CA", X"91", X"6F", X"01", X"79", X"75", X"35", X"F3", X"F9", X"C8", X"4F", X"E9", X"7C", X"8D", X"F0", X"16", X"DF", X"4B", X"BD", X"C8", X"5C", X"2C", X"EB", X"30", X"76", X"ED", X"E1", X"34", X"3E", X"98", X"F2", X"C2", X"BC", X"18", X"FA", X"94", X"7A", X"3D", X"5E", X"45", X"6E", X"FD", X"40", X"6C", X"A5", X"DF", X"8C", X"1C", X"0D", X"2F", X"F5", X"2A", X"31", X"A1", X"6D", X"7D", X"BD", X"6E", X"41", X"39", X"81", X"22", X"D0", X"16", X"2F", X"58", X"53", X"38", X"A3", X"C2", X"D2", X"2C", X"F0", X"5C", X"1C", X"4F", X"A6", X"D6", X"01", X"AC", X"19", X"D6", X"8D", X"31", X"D1", X"0B", X"27", X"97", X"81", X"9F", X"25", X"68", X"2C", X"FE", X"3F", X"75", X"25", X"B6", X"0E", X"01", X"FF", X"D6", X"42", X"EB", X"3B", X"5F", X"03", X"6A", X"90", X"60", X"D6", X"2E", X"CC", X"C6", X"54", X"DA", X"9C", X"69", X"1F", X"94", X"2D", X"41", X"6C", X"AF", X"66", X"A7", X"27", X"15", X"36", X"86", X"6F", X"4C", X"FF", X"5E", X"07", X"E7", X"D0", X"BD", X"8E", X"67", X"DC", X"53", X"BF", X"67", X"69", X"F8", X"38", X"88", X"FD", X"57", X"B2", X"EA", X"EC", X"BA", X"E5", X"2E", X"C1", X"6B", X"41", X"80", X"40", X"82", X"1D", X"A9", X"A6", X"58", X"FB", X"74", X"FE", X"58", X"67", X"EB", X"77", X"44", X"B8", X"84", X"58", X"BC", X"39", X"26", X"49", X"FE", X"1A", X"D7", X"DF", X"28", X"A7", X"4C", X"5A", X"9A", X"11", X"F0", X"5B", X"37", X"F0", X"C4", X"16", X"F3", X"08", X"7A", X"55", X"67", X"39", X"B5", X"D8", X"3A", X"A2", X"A5", X"FF", X"55", X"FB", X"71", X"D1", X"E4", X"F9", X"48", X"57", X"FA", X"5D", X"A8", X"7E", X"96", X"5B", X"1A", X"28", X"66", X"02", X"19", X"A2", X"CE", X"A4", X"BA", X"62", X"EC", X"41", X"7C", X"5C", X"E8", X"D6", X"67", X"5D", X"A2", X"B1", X"DC", X"78", X"C5", X"15", X"98", X"F9", X"DE", X"75", X"7A", X"E4", X"B6", X"84", X"95", X"47", X"A4", X"77", X"D4", X"94", X"D6", X"B4", X"CF", X"E7", X"29", X"24", X"31", X"E9", X"23", X"BF", X"CC", X"2B", X"BE", X"89", X"DB", X"DA", X"16", X"39", X"0A", X"0E", X"8A", X"43", X"F1", X"F6", X"49", X"F4", X"95", X"D0", X"48", X"5D", X"B1", X"DD", X"9A", X"FE", X"CB", X"65", X"7B", X"49", X"F9", X"4B", X"6C", X"AB", X"31", X"CD", X"B9", X"41", X"2B", X"FD", X"46", X"C5", X"0D", X"AB", X"16", X"8A", X"E6", X"BF", X"3F", X"F8", X"A9", X"D9", X"31", X"66", X"62", X"C2", X"0D", X"B7", X"66", X"88", X"9E", X"3F", X"DC", X"E6", X"C6", X"99", X"1D", X"3F", X"61", X"62", X"AA", X"F4", X"8F", X"4F", X"7B", X"FC", X"61", X"C7", X"04", X"2F", X"39", X"31", X"DA", X"87", X"FD", X"A0", X"B7", X"C4", X"DA", X"9C", X"E2", X"8F", X"6B", X"E2", X"EB", X"26", X"2B", X"04", X"4C", X"3E", X"A5", X"F1", X"D7", X"F9", X"CE", X"86", X"09", X"53", X"4D", X"E0", X"15", X"C3", X"F9", X"6F", X"E3", X"D9", X"DE", X"B3", X"C0", X"4B", X"F8", X"6D", X"89", X"B6", X"32", X"A3", X"70", X"98", X"E8", X"6D", X"19", X"8A", X"15", X"03", X"9D", X"CA", X"7E", X"66", X"F7", X"6B", X"1C", X"59", X"0B", X"A2", X"99", X"8B", X"03", X"DB", X"5C", X"83", X"09", X"7B", X"9B", X"6E", X"66", X"51", X"F8", X"87", X"CC", X"48", X"20", X"4F", X"E3", X"5B", X"A7", X"2D", X"03", X"A0", X"C8", X"EE", X"49", X"BE", X"7D", X"F9", X"8B", X"F3", X"6C", X"A8", X"C4", X"49", X"FA", X"08", X"2B", X"94", X"1A", X"A4", X"CA", X"D6", X"FD", X"AE", X"84", X"61", X"A0", X"70", X"E5", X"3C", X"4D", X"F3", X"8E", X"F1", X"E6", X"FD", X"8E", X"94", X"0F", X"0F", X"D0", X"89", X"C2", X"47", X"58", X"10", X"CA", X"BC", X"36", X"0B", X"D8", X"57", X"ED", X"43", X"39", X"C8", X"51", X"24", X"B2", X"76", X"F7", X"ED", X"1D", X"B4", X"01", X"08", X"CC", X"A9", X"8F", X"F6", X"3C", X"9D", X"77", X"31", X"AD", X"13", X"90", X"D3", X"81", X"51", X"F7", X"75", X"CC", X"4C", X"94", X"AC", X"A7", X"A0", X"36", X"7D", X"E1", X"8B", X"AC", X"63", X"1D", X"CC", X"48", X"78", X"25", X"4B", X"D6", X"40", X"DE", X"8F", X"36", X"54", X"9D", X"51", X"10", X"63", X"25", X"39", X"C3", X"49", X"7B", X"56", X"7A", X"D1", X"A7", X"23", X"7E", X"DC", X"47", X"E6", X"C1", X"98", X"A2", X"4D", X"C6", X"04", X"FE", X"AD", X"15", X"D6", X"93", X"99", X"79", X"7B", X"C6", X"61", X"5E", X"4D", X"33", X"0A", X"F2", X"25", X"CC", X"3C", X"A2", X"4A", X"F1", X"18", X"D3", X"A6", X"50", X"1C", X"62", X"92", X"0B", X"0A", X"B8", X"C5", X"43", X"1B", X"7A", X"EE", X"69", X"49", X"9D", X"C7", X"2F", X"3E", X"28", X"56", X"62", X"47", X"04", X"28", X"C1", X"75", X"C9", X"FA", X"B5", X"67", X"57", X"DD", X"9C", X"0B", X"F4", X"78", X"0D", X"47", X"22", X"B5", X"5B", X"59", X"20", X"76", X"23", X"93", X"91", X"FF", X"9E", X"A4", X"32", X"D2", X"2D", X"E0", X"5A", X"0F", X"C1", X"3E", X"AB", X"52", X"8E", X"DD", X"F3", X"FC", X"0C", X"97", X"0C", X"45", X"38", X"4A", X"C5", X"59", X"28", X"53", X"28", X"C9", X"1B", X"1D", X"97", X"EC", X"CD", X"EA", X"47", X"30", X"D2", X"9B", X"4A", X"E6", X"6A", X"81", X"1C", X"44", X"A0", X"58", X"BC", X"0C", X"93", X"41", X"1A", X"0E", X"49", X"34", X"90", X"60", X"8D", X"C1", X"EF", X"EA", X"B8", X"CA", X"D6", X"AB", X"E9", X"71", X"3B", X"7E", X"91", X"1A", X"0C", X"3A", X"1E", X"80", X"03", X"E3", X"92", X"11", X"3E", X"FA", X"97", X"65", X"7F", X"C7", X"62", X"D7", X"A2", X"4C", X"07", X"3F", X"7F", X"59", X"02", X"00", X"24", X"AB", X"E2", X"42", X"63", X"C6", X"C4", X"BA", X"B0", X"58", X"EE", X"1B", X"67", X"F3", X"EA", X"2F", X"4A", X"96", X"D0", X"F6", X"90", X"48", X"5B", X"51", X"78", X"90", X"87", X"0A", X"22", X"DC", X"C0", X"FA", X"90", X"06", X"05", X"32", X"A8", X"C0", X"F8", X"71", X"8F", X"EB", X"4D", X"AA", X"69", X"27", X"06", X"04", X"E6", X"CF", X"57", X"E6", X"BC", X"35", X"51", X"88", X"77", X"69", X"01", X"8E", X"0E", X"51", X"F2", X"2A", X"B2", X"21", X"4F", X"50", X"25", X"A8", X"B9", X"18", X"ED", X"E0", X"B5", X"20", X"CF", X"F3", X"62", X"DD", X"A9", X"8C", X"81", X"E1", X"3D", X"B0", X"9B", X"39", X"C6", X"00", X"45", X"7E", X"4B", X"98", X"95", X"80", X"54", X"5C", X"48", X"D2", X"36", X"C1", X"C8", X"F2", X"6A", X"F3", X"D8", X"7E", X"1A", X"70", X"8D", X"BE", X"56", X"7F", X"E1", X"E4", X"44", X"11", X"94", X"FA", X"AA", X"FF", X"40", X"32", X"FD", X"AA", X"46", X"27", X"68", X"7F", X"B7", X"BE", X"9F", X"49", X"E6", X"92", X"A6", X"51", X"08", X"A0", X"2E", X"38", X"03", X"DE", X"AB", X"18", X"FB", X"DC", X"99", X"5D", X"F0", X"6D", X"97", X"CC", X"B4", X"7B", X"40", X"1D", X"2F", X"5B", X"BB", X"44", X"41", X"AA", X"3F", X"B8", X"64", X"23", X"66", X"B8", X"07", X"4B", X"54", X"A0", X"A4", X"A2", X"C9", X"97", X"D7", X"9F", X"FF", X"27", X"91", X"F9", X"97", X"3B", X"EB", X"91", X"EF", X"C7", X"7B", X"C6", X"AF", X"95", X"B6", X"B9", X"01", X"F7", X"4C", X"B9", X"F9", X"DE", X"EA", X"F3", X"A1", X"66", X"D9", X"07", X"AC", X"40", X"42", X"2C", X"22", X"7F", X"CB", X"7C", X"AF", X"8C", X"F9", X"99", X"99", X"EF", X"D8", X"D9", X"99", X"14", X"EA", X"55", X"6A", X"D8", X"18", X"55", X"06", X"79", X"33", X"41", X"6C", X"8C", X"57", X"D9", X"CE", X"3C", X"AB", X"81", X"CF", X"26", X"80", X"1F", X"99", X"1C", X"FB", X"9C", X"1A", X"77", X"55", X"37", X"0C", X"4F", X"60", X"82", X"4F", X"B1", X"55", X"5C", X"B6", X"BE", X"61", X"F1", X"48", X"5B", X"93", X"6F", X"C3", X"95", X"82", X"1D", X"CD", X"23", X"D8", X"88", X"8B", X"71", X"A6", X"95", X"6D", X"79", X"BB", X"1B", X"92", X"AA", X"37", X"27", X"93", X"1B", X"EA", X"23", X"27", X"6B", X"C4", X"47", X"69", X"49", X"D9", X"16", X"B3", X"70", X"FF", X"F4", X"11", X"E0", X"DA", X"9C", X"6C", X"9C", X"CA", X"EF", X"60", X"37", X"8E", X"74", X"F5", X"77", X"CE", X"FB", X"FD", X"37", X"3E", X"1F", X"45", X"EF", X"FF", X"EE", X"8C", X"EF", X"EB", X"1F", X"84", X"D4", X"46", X"06", X"78", X"9A", X"07", X"68", X"08", X"4A", X"C0", X"51", X"92", X"14", X"6A", X"72", X"56", X"EE", X"91", X"82", X"2E", X"36", X"D6", X"F5", X"A5", X"80", X"22", X"20", X"80", X"42", X"4A", X"21", X"99", X"2E", X"E1", X"16", X"19", X"BC", X"08", X"98", X"D0", X"14", X"75", X"4F", X"B4", X"FD", X"4C", X"3C", X"EE", X"DC", X"66", X"52", X"AA", X"90", X"F9", X"4D", X"67", X"32", X"A1", X"F4", X"F4", X"41", X"26", X"3E", X"7C", X"BF", X"EC", X"48", X"23", X"52", X"40", X"FF", X"41", X"00", X"C1", X"F9", X"CD", X"C3", X"1F", X"B6", X"73", X"26", X"4B", X"2A", X"FC", X"B1", X"19", X"E1", X"DD", X"FE", X"C0", X"30", X"75", X"BF", X"75", X"2B", X"41", X"64", X"6C", X"70", X"73", X"75", X"02", X"83", X"1D", X"28", X"43", X"13", X"B8", X"32", X"16", X"C1", X"63", X"58", X"58", X"BA", X"CC", X"8E", X"41", X"28", X"02", X"50", X"B0", X"B5", X"30", X"DB", X"D6", X"6D", X"39", X"39", X"C8", X"DF", X"1A", X"5C", X"9A", X"08", X"49", X"9B", X"D1", X"62", X"1A", X"02", X"74", X"EC", X"DE", X"E7", X"59", X"8B", X"6F", X"1A", X"22", X"15", X"70", X"B3", X"CF", X"8E", X"8C", X"B7", X"02", X"25", X"76", X"70", X"7D");
signal frame_3: FRAME3 := (X"16", X"DC", X"C6", X"B4", X"09", X"09", X"B9", X"39", X"2B", X"07", X"08", X"86", X"C6", X"75", X"B1", X"04", X"23", X"E3", X"EB", X"C7", X"57", X"D0", X"77", X"63", X"02", X"EB", X"4A", X"A2", X"FD", X"99", X"1F", X"D0", X"47", X"EB", X"DA", X"45", X"6B", X"92", X"8F", X"A3", X"B9", X"88", X"29", X"8F", X"2C", X"5F", X"B8", X"AD", X"F7", X"E6", X"98", X"62", X"A5", X"C4", X"96", X"90", X"53", X"E4", X"D2", X"07", X"0C", X"86", X"0A", X"CE", X"6E", X"4C", X"25", X"61", X"86", X"67", X"D0", X"98", X"74", X"86", X"4E", X"1C", X"82", X"BB", X"23", X"B5", X"20", X"84", X"18", X"B8", X"17", X"8D", X"C7", X"46", X"3C", X"25", X"D2", X"C0", X"95", X"B0", X"17", X"DD", X"3C", X"4C", X"58", X"4B", X"9F", X"23", X"EE", X"E8", X"35", X"B0", X"93", X"EF", X"CD", X"7C", X"3A", X"AF", X"D7", X"F6", X"8A", X"2B", X"B6", X"DD", X"72", X"97", X"71", X"77", X"12", X"B8", X"3A", X"F2", X"63", X"7A", X"DC", X"C3", X"70", X"89", X"F1", X"81", X"21", X"96", X"84", X"44", X"7D", X"1B", X"FF", X"E4", X"F4", X"AC", X"19", X"52", X"02", X"4C", X"DE", X"21", X"D6", X"F1", X"21", X"6B", X"FF", X"97", X"B1", X"A1", X"B9", X"1C", X"1E", X"AD", X"7F", X"A3", X"BD", X"5A", X"3B", X"FF", X"02", X"FC", X"D0", X"2A", X"49", X"2A", X"35", X"C9", X"F4", X"FF", X"6A", X"99", X"26", X"EF", X"8A", X"9C", X"7B", X"99", X"00", X"E2", X"09", X"32", X"94", X"27", X"7B", X"6C", X"2F", X"00", X"33", X"39", X"52", X"51", X"0C", X"3B", X"24", X"D1", X"BC", X"D7", X"EB", X"91", X"EE", X"B9", X"4D", X"F1", X"B8", X"23", X"B9", X"E1", X"4F", X"47", X"B7", X"D0", X"2B", X"EF", X"C0", X"83", X"2B", X"B7", X"00", X"3B", X"D0", X"1F", X"06", X"34", X"47", X"FD", X"80", X"92", X"7A", X"F2", X"DC", X"E2", X"C2", X"33", X"52", X"BB", X"CC", X"F8", X"E6", X"89", X"E9", X"5C", X"ED", X"F9", X"01", X"7B", X"0F", X"76", X"6A", X"B8", X"42", X"3B", X"8F", X"E9", X"9B", X"7F", X"5B", X"D5", X"FF", X"AE", X"FF", X"96", X"A0", X"A5", X"5C", X"4E", X"14", X"A1", X"57", X"D8", X"71", X"F7", X"9D", X"8C", X"A8", X"16", X"F1", X"24", X"57", X"26", X"EA", X"66", X"D7", X"C1", X"77", X"E3", X"9F", X"15", X"1E", X"BA", X"5E", X"90", X"F3", X"0B", X"55", X"9C", X"F2", X"3B", X"38", X"33", X"6E", X"36", X"0C", X"CF", X"BB", X"AF", X"E3", X"D1", X"BB", X"1A", X"D6", X"C5", X"35", X"12", X"95", X"03", X"A1", X"2B", X"82", X"92", X"B4", X"E0", X"4E", X"AA", X"F0", X"47", X"91", X"74", X"D1", X"A4", X"FF", X"90", X"F7", X"0C", X"7E", X"68", X"B7", X"FF", X"CD", X"18", X"74", X"FE", X"41", X"34", X"A0", X"10", X"6D", X"D5", X"5B", X"20", X"E0", X"66", X"60", X"58", X"47", X"71", X"8D", X"CA", X"2F", X"D3", X"D2", X"DA", X"2A", X"90", X"6E", X"76", X"6C", X"53", X"FE", X"6E", X"7D", X"A4", X"56", X"60", X"75", X"50", X"4F", X"F1", X"A8", X"71", X"27", X"21", X"57", X"A5", X"D1", X"42", X"2F", X"1E", X"FE", X"CD", X"1F", X"6B", X"31", X"65", X"30", X"B3", X"D1", X"4F", X"B7", X"A9", X"85", X"5E", X"8E", X"D4", X"BE", X"AB", X"F4", X"43", X"ED", X"C4", X"AE", X"8B", X"8E", X"1F", X"AB", X"85", X"D4", X"C3", X"C4", X"29", X"B9", X"2B", X"95", X"87", X"FE", X"A5", X"F2", X"7A", X"7D", X"61", X"B9", X"B9", X"CC", X"1B", X"92", X"C4", X"BB", X"AC", X"15", X"B6", X"65", X"FB", X"16", X"61", X"3F", X"6E", X"DD", X"AC", X"DA", X"52", X"11", X"D8", X"92", X"7A", X"8B", X"74", X"7E", X"B1", X"5C", X"10", X"49", X"3F", X"09", X"66", X"6A", X"97", X"BC", X"4C", X"D9", X"63", X"28", X"FD", X"1B", X"42", X"C3", X"03", X"2D", X"D2", X"76", X"5F", X"53", X"59", X"56", X"87", X"0C", X"0F", X"5C", X"F6", X"4B", X"DB", X"2E", X"74", X"B3", X"D1", X"39", X"BA", X"0D", X"1A", X"63", X"DB", X"60", X"27", X"A7", X"44", X"C4", X"EB", X"4D", X"E6", X"D6", X"7F", X"6D", X"CA", X"08", X"BF", X"06", X"37", X"0A", X"8E", X"B4", X"00", X"A9", X"07", X"66", X"8A", X"DD", X"AA", X"05", X"B2", X"31", X"51", X"88", X"43", X"F2", X"06", X"90", X"E4", X"FF", X"7B", X"8F", X"CC", X"F5", X"E3", X"2C", X"F2", X"11", X"61", X"18", X"5A", X"B7", X"B5", X"FE", X"15", X"E7", X"53", X"04", X"C4", X"32", X"A4", X"79", X"39", X"E8", X"96", X"C2", X"E1", X"82", X"67", X"1F", X"6D", X"9E", X"1D", X"64", X"FA", X"34", X"4A", X"34", X"8E", X"44", X"9D", X"2C", X"78", X"D3", X"53", X"10", X"7B", X"30", X"8E", X"08", X"A2", X"2B", X"F7", X"A7", X"37", X"8D", X"7B", X"92", X"78", X"2B", X"DE", X"38", X"44", X"2D", X"A1", X"C9", X"10", X"05", X"82", X"CF", X"87", X"10", X"7C", X"DD", X"22", X"20", X"9C", X"7C", X"C9", X"46", X"DA", X"75", X"AA", X"5E", X"B2", X"71", X"60", X"58", X"79", X"4A", X"AD", X"6B", X"35", X"2E", X"30", X"89", X"04", X"58", X"B6", X"0A", X"D0", X"E0", X"94", X"77", X"09", X"CD", X"52", X"75", X"65", X"FF", X"D9", X"6F", X"4F", X"96", X"AE", X"5A", X"C2", X"BA", X"7A", X"BD", X"84", X"7F", X"4B", X"03", X"2C", X"02", X"42", X"E6", X"DB", X"C5", X"8D", X"98", X"ED", X"91", X"56", X"D2", X"46", X"94", X"0B", X"94", X"E5", X"84", X"A4", X"B6", X"8F", X"35", X"47", X"9A", X"70", X"DA", X"3E", X"65", X"8D", X"99", X"AD", X"F9", X"CD", X"F4", X"D7", X"DA", X"F7", X"D1", X"D2", X"72", X"02", X"D9", X"02", X"2F", X"67", X"0A", X"31", X"97", X"7E", X"49", X"6B", X"8D", X"8C", X"A3", X"8A", X"19", X"2B", X"4F", X"7F", X"B8", X"BC", X"AA", X"EB", X"02", X"0F", X"F7", X"40", X"18", X"C2", X"61", X"57", X"25", X"D7", X"86", X"61", X"C6", X"7E", X"F1", X"AF", X"C9", X"5D", X"FD", X"7E", X"77", X"7F", X"D7", X"C2", X"7E", X"E5", X"C0", X"57", X"10", X"6C", X"94", X"1B", X"DB", X"EC", X"91", X"1C", X"73", X"94", X"9B", X"9D", X"31", X"74", X"E8", X"B7", X"5B", X"14", X"C1", X"BA", X"D2", X"E5", X"07", X"B8", X"37", X"D1", X"4A", X"66", X"1B", X"EB", X"5E", X"BD", X"42", X"A3", X"13", X"D5", X"C9", X"9A", X"82", X"26", X"45", X"C7", X"6B", X"E1", X"E5", X"5B", X"8C", X"66", X"60", X"77", X"A2", X"40", X"D8", X"9F", X"C8", X"14", X"E9", X"53", X"4B", X"C8", X"52", X"C1", X"77", X"90", X"04", X"7C", X"1F", X"25", X"F7", X"6D", X"4B", X"00", X"74", X"27", X"E0", X"E0", X"26", X"DD", X"BE", X"67", X"DE", X"7F", X"17", X"D7", X"FA", X"5E", X"D0", X"DB", X"00", X"E2", X"A8", X"A1", X"36", X"3B", X"29", X"71", X"E8", X"97", X"E7", X"03", X"45", X"E3", X"31", X"BF", X"A3", X"34", X"12", X"ED", X"48", X"C3", X"B2", X"1B", X"98", X"36", X"FE", X"36", X"63", X"95", X"17", X"F7", X"B3", X"98", X"49", X"20", X"C6", X"42", X"FB", X"3D", X"0F", X"20", X"86", X"CF", X"A3", X"66", X"39", X"19", X"D7", X"A2", X"12", X"C4", X"1F", X"88", X"B9", X"0A", X"CB", X"0C", X"53", X"B4", X"8E", X"A8", X"E2", X"9F", X"94", X"3A", X"BB", X"58", X"3C", X"B8", X"74", X"25", X"2C", X"E7", X"B5", X"22", X"99", X"C0", X"A4", X"5B", X"06", X"5B", X"58", X"00", X"C8", X"ED", X"5B", X"5F", X"03", X"BB", X"C8", X"AD", X"BF", X"10", X"06", X"E4", X"FD", X"FC", X"E0", X"1C", X"B8", X"2A", X"0A", X"76", X"2C", X"7E", X"E4", X"05", X"07", X"B4", X"8D", X"C4", X"58", X"EF", X"2B", X"1E", X"EC", X"C9", X"E1", X"CA", X"29", X"C9", X"C2", X"4C", X"0F", X"DA", X"44", X"72", X"0A", X"44", X"BB", X"B2", X"F4", X"8D", X"06", X"24", X"3E", X"24", X"79", X"C9", X"02", X"85", X"1A", X"FE", X"86", X"7F", X"40", X"02", X"6A", X"83", X"8D", X"97", X"A7", X"F1", X"E3", X"52", X"44", X"52", X"B5", X"60", X"4A", X"DB", X"66", X"C5", X"34", X"81", X"E8", X"F9", X"DF", X"52", X"03", X"D9", X"08", X"C8", X"41", X"10", X"EE", X"1B", X"C7", X"F2", X"95", X"28", X"8C", X"FB", X"E9", X"90", X"DA", X"C9", X"7E", X"C6", X"2D", X"80", X"E8", X"BC", X"3B", X"95", X"A4", X"CE", X"A1", X"6F", X"C2", X"97", X"94", X"3D", X"C4", X"3E", X"B3", X"B4", X"58", X"84", X"2E", X"7C", X"FD", X"F8", X"83", X"D1", X"CD", X"A9", X"D8", X"E8", X"D1", X"0F", X"0E", X"36", X"6F", X"4C", X"55", X"01", X"CD", X"14", X"A6", X"91", X"20", X"43", X"E5", X"32", X"C9", X"BE", X"97", X"EB", X"7D", X"55", X"76", X"4F", X"DD", X"03", X"3F", X"0B", X"03", X"17", X"83", X"36", X"FA", X"B2", X"97", X"95", X"D5", X"14", X"57", X"BA", X"68", X"1B", X"E1", X"24", X"64", X"41", X"71", X"5A", X"FB", X"C4", X"88", X"33", X"73", X"92", X"75", X"61", X"67", X"59", X"8D", X"BE", X"89", X"2E", X"5E", X"97", X"50", X"85", X"04", X"EA", X"F2", X"A9", X"1D", X"C7", X"3F", X"5F", X"65", X"A1", X"A9", X"D8", X"39", X"2C", X"F8", X"E8", X"46", X"94", X"F6", X"D4", X"30", X"4D", X"43", X"55", X"47", X"21", X"A7", X"10", X"A4", X"05", X"E4", X"FB", X"B3", X"22", X"E9", X"62", X"10", X"7D", X"7E", X"8C", X"76", X"B5", X"44", X"A5", X"AD", X"3D", X"5C", X"3E", X"5A", X"15", X"33", X"C2", X"83", X"DC", X"FB", X"C6", X"F6", X"B6", X"A5", X"C5", X"C5", X"16", X"77", X"E5", X"96", X"1B", X"09", X"60", X"AB", X"CA", X"E1", X"A1", X"51", X"DF", X"F3", X"A2", X"AB", X"8F", X"D6", X"57", X"74", X"E7", X"3D", X"DE", X"CE", X"BD", X"45", X"34", X"EF", X"50", X"BB", X"82", X"27", X"6A", X"84", X"4D", X"2E", X"CD", X"C5", X"6C", X"79", X"73", X"EE", X"7C", X"78", X"11", X"A1", X"77", X"57", X"4F", X"58", X"B5", X"C0", X"A2", X"6C", X"64", X"F6", X"B0", X"7D", X"8B", X"A3", X"7C", X"C8", X"D1", X"CD", X"1C", X"E2", X"9F", X"7B", X"9B", X"12", X"D2", X"A2", X"50", X"75", X"75", X"C6", X"4A", X"31", X"33", X"20", X"B7", X"B2", X"69", X"5B", X"DA", X"82", X"5E", X"44", X"C1", X"73", X"50", X"88", X"BD", X"B5", X"1B", X"69", X"FC", X"CB", X"0F", X"13", X"30", X"2E", X"70", X"D3", X"2A", X"94", X"0F", X"48", X"8F", X"ED", X"79", X"1C", X"9D", X"A3", X"BC", X"40", X"FF", X"DB", X"85", X"7D", X"0A", X"1A", X"84", X"13", X"8A", X"AC", X"E7", X"5C", X"51", X"AB", X"B9", X"11", X"94", X"2B", X"14", X"34", X"D9", X"69", X"F8", X"F5", X"5C", X"3F", X"17", X"C3", X"42", X"8B", X"3B", X"33", X"34", X"12", X"97", X"6E", X"F8", X"8D", X"A0", X"0D", X"55", X"1C", X"BA", X"DF", X"F2", X"42", X"14", X"65", X"D5", X"D3", X"6F", X"57", X"85", X"70", X"C7", X"C6", X"12", X"E9", X"65", X"45", X"1A", X"9C", X"1E", X"44", X"9D", X"AE", X"D0", X"85", X"8D", X"0E", X"42", X"52", X"31", X"53", X"4B", X"E7", X"54", X"85", X"17", X"60", X"04", X"10", X"B7", X"58", X"F7", X"60", X"62", X"73", X"04", X"51");

begin

o_src_ip <=  x"f0000000"; 
o_dst_ip <=  x"00000002"; 
o_src_port <= x"0f00";
o_dst_port <= x"0002";
o_active_mode <= '1';
o_timeout <= (others => '1');


stim1: process(clk, reset)
begin
  tx_tlast <= '0';
  if(rising_edge(clk) and reset = '1') then
    i <= 0;
	state <= start_trans;
  elsif (rising_edge(clk)) then
    case state is
	  when start_trans =>
	    o_start <= '1';
		o_open <= '1';
	    if (i_close = '1') then
			state <= send_frame1;
		end if;
	  when send_frame1 =>
	   tx_tvalid <= '1';
	   tx_tdata  <= frame_1(i);
	   if(tx_tready = '1') then
	     i <= i + 1;
	     if(i = 50) then
	       state <= send_frame2;
		   tx_tlast <= '1';
		   i <= 0;
	     end if;
	   end if;
	  when send_frame2 =>
	    tx_tvalid <= '1';
		tx_tdata <= frame_2(i);
		if(tx_tready = '1') then
		  i <= i + 1;
		  if(i = 4200) then
		    state <= send_frame3;
		    tx_tlast <= '1';
			i <= 0;
		  end if;
		end if;
	  when send_frame3 =>
	    tx_tvalid <= '1';
		tx_tdata <= frame_3(i);
		if(tx_tready = '1') then
		  i <= i + 1;
		  if(i = 1400) then
		    state <= request_close;
		    tx_tlast <= '1';
		  end if;
		end if;
	  when request_close =>
	    o_open <= '0';
	end case;
  end if;
end process;
end behavioural;